/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none 
 
module tt_um_uwasic_dinogame (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);


  wire [8:0] obstacle1_pos;
  wire [8:0] obstacle2_pos;
  wire [2:0] obstacle1_type;
  wire [2:0] obstacle2_type;
  wire [7:0] rng;
  wire gametick;
  obstacles #(.GEN_LINE(250)) obstacles_inst (
      .clk(gametick),
      .rst_n(rst_n),
      .rng(rng),
      .obstacle1_pos(obstacle1_pos),
      .obstacle2_pos(obstacle2_pos),
      .obstacle1_type(obstacle1_type),
      .obstacle2_type(obstacle2_type)
  );


  // All output pins must be assigned. If not used, assign to 0.
  assign uo_out  = ui_in + uio_in;  // Example: ou_out is the sum of ui_in and uio_in
  assign uio_out = 0;
  assign uio_oe  = 0;

  // List all unused inputs to prevent warnings
  wire _unused = &{ena, clk, rst_n, 1'b0};

endmodule
